//from Cello UCF Supplemental

module x01(output out, input a, b, c);
    and(out, a, b, c); 
endmodule