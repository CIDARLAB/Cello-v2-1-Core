module Main(in1, out1);
  output out1;
  input in1;  
  
  assign g1 = ~in1;
  
  assign out1 = g1;
  
  endmodule
  
 // Single Not Gate
 // Total Gates: 3
 // Gates: 1, 40, 52
